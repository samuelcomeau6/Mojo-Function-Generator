module transmit_rom (
    input clk,
    input [7:0] mess,
    input [3:0] addr,
    output [7:0] data
  );
 
  wire [7:0] rom_data [13:0][17:0];
 
  assign rom_data[0][1] = " ";
  assign rom_data[1][1] = "S";
  assign rom_data[2][1] = "q";
  assign rom_data[3][1] = "u";
  assign rom_data[4][1] = "a";
  assign rom_data[5][1] = "r";
  assign rom_data[6][1] = "e";
  assign rom_data[7][1] = " ";
  assign rom_data[8][1] = "W";
  assign rom_data[9][1] = "a";
  assign rom_data[10][1] = "v";
  assign rom_data[11][1] = "e";
  assign rom_data[12][1] = "\n";
  assign rom_data[13][1] = "\r";
  assign rom_data[0][2] = " ";
  assign rom_data[1][2] = "S";
  assign rom_data[2][2] = "i";
  assign rom_data[3][2] = "n";
  assign rom_data[4][2] = "e";
  assign rom_data[5][2] = " ";
  assign rom_data[6][2] = "W";
  assign rom_data[7][2] = "a";
  assign rom_data[8][2] = "v";
  assign rom_data[9][2] = "e";
  assign rom_data[10][2] = " ";
  assign rom_data[11][2] = " ";
  assign rom_data[12][2] = "\n";
  assign rom_data[13][2] = "\r";
  assign rom_data[0][3]= " ";
  assign rom_data[1][3] = "T";
  assign rom_data[2][3] = "r";
  assign rom_data[3][3] = "i";
  assign rom_data[4][3] = " ";
  assign rom_data[5][3] = "W";
  assign rom_data[6][3] = "a";
  assign rom_data[7][3] = "v";
  assign rom_data[8][3] = "e";
  assign rom_data[9][3] = " ";
  assign rom_data[10][3] = " ";
  assign rom_data[11][3] = " ";
  assign rom_data[12][3] = "\n";
  assign rom_data[13][3] = "\r"; 
  assign rom_data[0][4] = " ";
  assign rom_data[1][4] = "S";
  assign rom_data[2][4] = "a";
  assign rom_data[3][4] = "w";
  assign rom_data[4][4] = " ";
  assign rom_data[5][4] = "W";
  assign rom_data[6][4] = "a";
  assign rom_data[7][4] = "v";
  assign rom_data[8][4] = "e";
  assign rom_data[9][4] = " ";
  assign rom_data[10][4] = " ";
  assign rom_data[11][4] = " ";
  assign rom_data[12][4] = "\n";
  assign rom_data[13][4] = "\r"; 
  assign rom_data[0][5] = " ";
  assign rom_data[1][5] = "R";
  assign rom_data[2][5] = "a";
  assign rom_data[3][5] = "i";
  assign rom_data[4][5] = "s";
  assign rom_data[5][5] = "e";
  assign rom_data[6][5] = " ";
  assign rom_data[7][5] = "F";
  assign rom_data[8][5] = "r";
  assign rom_data[9][5] = "e";
  assign rom_data[10][5] = "q";
  assign rom_data[11][5] = " ";
  assign rom_data[12][5] = "\n";
  assign rom_data[13][5] = "\r"; 
  assign rom_data[0][6] = " ";
  assign rom_data[1][6] = "L";
  assign rom_data[2][6] = "o";
  assign rom_data[3][6] = "w";
  assign rom_data[4][6] = "e";
  assign rom_data[5][6] = "r";
  assign rom_data[6][6] = " ";
  assign rom_data[7][6] = "F";
  assign rom_data[8][6] = "r";
  assign rom_data[9][6] = "e";
  assign rom_data[10][6] = "q";
  assign rom_data[11][6] = " ";
  assign rom_data[12][6] = "\n";
  assign rom_data[13][6] = "\r"; 
  assign rom_data[0][7] = " ";
  assign rom_data[1][7] = "R";
  assign rom_data[2][7] = "s";
  assign rom_data[3][7] = "t";
  assign rom_data[4][7] = " ";
  assign rom_data[5][7] = "f";
  assign rom_data[6][7] = "=";
  assign rom_data[7][7] = "2";
  assign rom_data[8][7] = "k";
  assign rom_data[9][7] = "H";
  assign rom_data[10][7] = "a";
  assign rom_data[11][7] = " ";
  assign rom_data[12][7] = "\n";
  assign rom_data[13][7] = "\r"; 
  assign rom_data[0][8] = " ";
  assign rom_data[1][8] = "S";
  assign rom_data[2][8] = "e";
  assign rom_data[3][8] = "t";
  assign rom_data[4][8] = " ";
  assign rom_data[5][8] = "f";
  assign rom_data[6][8] = "=";
  assign rom_data[7][8] = "1";
  assign rom_data[8][8] = "H";
  assign rom_data[9][8] = "z";
  assign rom_data[10][8] = " ";
  assign rom_data[11][8] = " ";
  assign rom_data[12][8] = "\n";
  assign rom_data[13][8] = "\r";
  assign rom_data[0][9] = " ";
  assign rom_data[1][9] = "S";
  assign rom_data[2][9] = "e";
  assign rom_data[3][9] = "t";
  assign rom_data[4][9] = " ";
  assign rom_data[5][9] = "f";
  assign rom_data[6][9] = "=";
  assign rom_data[7][9] = "1";
  assign rom_data[8][9] = "0";
  assign rom_data[9][9] = "H";
  assign rom_data[10][9] = "z";
  assign rom_data[11][9] = " ";
  assign rom_data[12][9] = "\n";
  assign rom_data[13][9] = "\r";  
  assign rom_data[0][10] = " ";
  assign rom_data[1][10] = "S";
  assign rom_data[2][10] = "e";
  assign rom_data[3][10] = "t";
  assign rom_data[4][10] = " ";
  assign rom_data[5][10] = "f";
  assign rom_data[6][10] = "=";
  assign rom_data[7][10] = "1";
  assign rom_data[8][10] = "0";
  assign rom_data[9][10] = "0";
  assign rom_data[10][10] = "H";
  assign rom_data[11][10] = "z";
  assign rom_data[12][10] = "\n";
  assign rom_data[13][10] = "\r"; 
  assign rom_data[0][11] = " ";
  assign rom_data[1][11] = "S";
  assign rom_data[2][11] = "e";
  assign rom_data[3][11] = "t";
  assign rom_data[4][11] = " ";
  assign rom_data[5][11] = "f";
  assign rom_data[6][11] = "=";
  assign rom_data[7][11] = "1";
  assign rom_data[8][11] = "k";
  assign rom_data[9][11] = "H";
  assign rom_data[10][11] = "z";
  assign rom_data[11][11] = " ";
  assign rom_data[12][11] = "\n";
  assign rom_data[13][11] = "\r";
  assign rom_data[0][12] = " ";
  assign rom_data[1][12] = "S";
  assign rom_data[2][12] = "e";
  assign rom_data[3][12] = "t";
  assign rom_data[4][12] = " ";
  assign rom_data[5][12] = "f";
  assign rom_data[6][12] = "=";
  assign rom_data[7][12] = "1";
  assign rom_data[8][12] = "0";
  assign rom_data[9][12] = "k";
  assign rom_data[10][12] = "H";
  assign rom_data[11][12] = "z";
  assign rom_data[12][12] = "\n";
  assign rom_data[13][12] = "\r";
  assign rom_data[0][13] = " ";
  assign rom_data[1][13] = "S";
  assign rom_data[2][13] = "e";
  assign rom_data[3][13] = "t";
  assign rom_data[4][13] = "f";
  assign rom_data[5][13] = "=";
  assign rom_data[6][13] = "1";
  assign rom_data[7][13] = "0";
  assign rom_data[8][13] = "0";
  assign rom_data[9][13] = "k";
  assign rom_data[10][13] = "H";
  assign rom_data[11][13] = "z";
  assign rom_data[12][13] = "\n";
  assign rom_data[13][13] = "\r";
  assign rom_data[0][14] = " ";
  assign rom_data[1][14] = "S";
  assign rom_data[2][14] = "e";
  assign rom_data[3][14] = "t";
  assign rom_data[4][14] = " ";
  assign rom_data[5][14] = "f";
  assign rom_data[6][14] = "=";
  assign rom_data[7][14] = "1";
  assign rom_data[8][14] = "M";
  assign rom_data[9][14] = "H";
  assign rom_data[10][14] = "z";
  assign rom_data[11][14] = " ";
  assign rom_data[12][14] = "\n";
  assign rom_data[13][14] = "\r";
  assign rom_data[0][15] = " ";
  assign rom_data[1][15] = "S";
  assign rom_data[2][15] = "e";
  assign rom_data[3][15] = "t";
  assign rom_data[4][15] = " ";
  assign rom_data[5][15] = "f";
  assign rom_data[6][15] = "=";
  assign rom_data[7][15] = "1";
  assign rom_data[8][15] = "0";
  assign rom_data[9][15] = "M";
  assign rom_data[10][15] = "H";
  assign rom_data[11][15] = "z";
  assign rom_data[12][15] = "\n";
  assign rom_data[13][15] = "\r";
  assign rom_data[0][16] = " ";
  assign rom_data[1][16] = "D";
  assign rom_data[2][16] = "o";
  assign rom_data[3][16] = "u";
  assign rom_data[4][16] = "b";
  assign rom_data[5][16] = "l";
  assign rom_data[6][16] = "e";
  assign rom_data[7][16] = " ";
  assign rom_data[8][16] = "F";
  assign rom_data[9][16] = "r";
  assign rom_data[10][16] = "e";
  assign rom_data[11][16] = "q";
  assign rom_data[12][16] = "\n";
  assign rom_data[13][16] = "\r";
  assign rom_data[0][17] = " ";
  assign rom_data[1][17] = "H";
  assign rom_data[2][17] = "a";
  assign rom_data[3][17] = "l";
  assign rom_data[4][17] = "f";
  assign rom_data[5][17] = " ";
  assign rom_data[6][17] = "F";
  assign rom_data[7][17] = "r";
  assign rom_data[8][17] = "e";
  assign rom_data[9][17] = "q";
  assign rom_data[10][17] = " ";
  assign rom_data[11][17] = " ";
  assign rom_data[12][17] = "\n";
  assign rom_data[13][17] = "\r";
    reg [7:0] data_d, data_q;
 
  assign data = data_q;
 
  always @(*) begin
    if (addr > 4'd13)
      data_d = " ";
    else
      data_d = rom_data[addr][mess];
  end
 
  always @(posedge clk) begin
    data_q <= data_d;
  end
 
endmodule
